
module display(diff, sinal, A, B, C, D, E, F, G, DP);
	
	input [3:0] diff;
	input sinal;
	output A, B, C, D, E, F, G, DP;

	
	wire SINAL_AND_NOT_DIFF2, DIFF2_AND_NOT_DIFF1_AND_NOT_DIFF0, DIFF2_AND_DIFF1_AND_DIFF0, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, NOT_DIFF_2_AND_NOT_DIFF1_AND_DIFF0, DIFF2_AND_NOT_DIFF0, DIFF1_AND_NOT_DIFF0, SINAL_AND_NOT_DIFF3, SINAL_AND_NOT_DIFF1, NOT_SINAL_AND_DIFF2, DIFF3_AND_NOT_DIFF2, NOT_DIFF1_AND_NOT_DIFF0, NOT_DIFF2_AND_NOT_DIFF1, DIFF2_AND_DIFF1_DIFF0;

	wire NOT_DIFF0, NOT_DIFF1, NOT_DIFF2, NOT_DIFF3, NOT_SINAL;
	not not0(NOT_DIFF0, diff[0]);
	not not1(NOT_DIFF1, diff[1]);
	not not2(NOT_DIFF2, diff[2]);
	not not3(NOT_DIFF3, diff[3]);
	not not4(NOT_SINAL, sinal);

	// Segmento A
	and andA0 (SINAL_AND_NOT_DIFF2, sinal, NOT_DIFF2);
	and andA1 (NOT_SINAL_AND_DIFF3, NOT_SINAL, diff[3]);
	and andA2 (NOT_DIFF3_AND_DIFF2, NOT_DIFF3, diff[2]);
	and andA3 (DIFF2_AND_DIFF1_DIFF0, diff[2], diff[1], diff[0]);
	and andA4 (DIFF2_AND_NOT_DIFF1_AND_NOT_DIFF0, diff[2], NOT_DIFF1, NOT_DIFF0);
	and andA5 (NOT_DIFF_2_AND_NOT_DIFF1_AND_DIFF0, NOT_DIFF2, NOT_DIFF1, diff[0]);

	or orA0 (A, SINAL_AND_NOT_DIFF2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, DIFF2_AND_DIFF1_DIFF0, DIFF2_AND_NOT_DIFF1_AND_NOT_DIFF0, NOT_DIFF_2_AND_NOT_DIFF1_AND_DIFF0);


	// Segmento B
	or orB0 (B, SINAL_AND_NOT_DIFF2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, DIFF2_AND_NOT_DIFF1_AND_NOT_DIFF0);

	// Segmento C
	and andC3 (DIFF2_AND_NOT_DIFF0, diff[2], NOT_DIFF0);
	and andC4 (DIFF1_AND_NOT_DIFF0, diff[1], NOT_DIFF0);

	or orC0 (C, SINAL_AND_NOT_DIFF2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, DIFF2_AND_NOT_DIFF0, DIFF1_AND_NOT_DIFF0);

	// Segmento D
	and andD0 (DIFF2_AND_DIFF1_AND_DIFF0, diff[2], diff[1], diff[0]);
	or orD0 (D, SINAL_AND_NOT_DIFF2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, DIFF2_AND_DIFF1_AND_DIFF0, DIFF2_AND_NOT_DIFF1_AND_NOT_DIFF0, NOT_DIFF_2_AND_NOT_DIFF1_AND_DIFF0);

	// Segmento E
	and andE0 (SINAL_AND_NOT_DIFF3, sinal, NOT_DIFF3);
	and andE1 (SINAL_AND_NOT_DIFF1, sinal, NOT_DIFF1);
	and andE2 (NOT_SINAL_AND_DIFF2, NOT_SINAL, diff[2]);
	and andE3 (DIFF3_AND_NOT_DIFF2, diff[3], NOT_DIFF2);

	or orE0 (E, SINAL_AND_NOT_DIFF3, SINAL_AND_NOT_DIFF1, NOT_SINAL_AND_DIFF2, DIFF3_AND_NOT_DIFF2, diff[0]);
	
	// Segmento F	
	or orF0 (F, sinal, diff[3], diff[2], diff[1], diff[0]);

	// Segmento G

	and andG1 (NOT_DIFF1_AND_NOT_DIFF0, NOT_DIFF1, NOT_DIFF0);
	and andG2 (NOT_DIFF2_AND_NOT_DIFF1, NOT_DIFF2, NOT_DIFF1);
	
	or orG0 (G, SINAL_AND_NOT_DIFF2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, DIFF2_AND_DIFF1_AND_DIFF0, NOT_DIFF2_AND_NOT_DIFF1, NOT_DIFF1_AND_NOT_DIFF0);
	

	// 	 A 			B			 C			D			E
	// sinal	diff3	 diff2	diff1	diff0

	// Segmento DP
	or orDP0 (DP, NOT_SINAL, NOT_DIFF3, NOT_DIFF2, NOT_DIFF1_AND_NOT_DIFF0);
	
endmodule 