
module display(diff, sinal, A, B, C, D, E, F, G, DP);
	
	input [3:0] diff;
	input sinal;
	output A, B, C, D, E, F, G, DP;
	
	wire SINAL_AND_NOT_DIFF_2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, NOT_DIFF0_AND_DIFF2, NOT_DIFF_2_AND_NOT_DIFF1_AND_DIFF0, DIFF2_AND_NOT_DIFF1_AND_NOT_DIFF0;
	wire DIFF2_AND_NOT_DIFF1, NOT_DIFF2_AND_DIFF1_AND_NOT_DIFF0, DIFF2_AND_NOT_DIFF0, NOT_DIFF2_AND_NOT_DIFF1_AND_DIFF_0,  SINAL_AND_NOT_DIFF_0, NOT_SINAL_AND_DIFF2, NOT_DIFF2_AND_DIFF0;	
	wire NOT_DIFF3_AND_DIFF1, SINAL_AND_DIFF1;
	
	wire NOT_DIFF0, NOT_DIFF1, NOT_DIFF2, NOT_DIFF3, NOT_SINAL;
	not not0(NOT_DIFF0, diff[0]);
	not not1(NOT_DIFF1, diff[1]);
	not not2(NOT_DIFF2, diff[2]);
	not not3(NOT_DIFF3, diff[3]);
	not not4(NOT_SINAL, sinal);
	
	// Segmento A
	and and0 (SINAL_AND_NOT_DIFF_2, sinal, NOT_DIFF2);
	and and1 (NOT_SINAL_AND_DIFF3, NOT_SINAL, diff[3]);
	and and2 (NOT_DIFF3_AND_DIFF2, NOT_DIFF3, diff[2]);
	and and3 (NOT_DIFF0_AND_DIFF2, NOT_DIFF0, diff[2]);
	and and4 (NOT_DIFF_2_AND_NOT_DIFF1_AND_DIFF0, NOT_DIFF2, NOT_DIFF1, diff[0]);
	or or0 (A, SINAL_AND_NOT_DIFF_2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, NOT_DIFF0_AND_DIFF2, NOT_DIFF_2_AND_NOT_DIFF1_AND_DIFF0);
	
	// Segmento B
	and and5 (DIFF2_AND_NOT_DIFF1_AND_NOT_DIFF0, diff[2], NOT_DIFF1, NOT_DIFF0);
	or or1 (B, SINAL_AND_NOT_DIFF_2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, DIFF2_AND_NOT_DIFF1_AND_NOT_DIFF0);
	
	// Segmento C
	and and6 (DIFF2_AND_NOT_DIFF1, diff[2], NOT_DIFF1);
	and and7 (NOT_DIFF2_AND_DIFF1_AND_NOT_DIFF0, NOT_DIFF2, diff[1], NOT_DIFF0);
	or or2 (C, SINAL_AND_NOT_DIFF_2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, DIFF2_AND_NOT_DIFF1, NOT_DIFF2_AND_DIFF1_AND_NOT_DIFF0);
	
	// Segmento D
	and and8 (DIFF2_AND_NOT_DIFF0, diff[2], NOT_DIFF0);
	and and9(NOT_DIFF2_AND_NOT_DIFF1_AND_DIFF_0, NOT_DIFF2, NOT_DIFF1, diff[0]);
	or or3 (D, SINAL_AND_NOT_DIFF_2, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, DIFF2_AND_NOT_DIFF0, NOT_DIFF2_AND_NOT_DIFF1_AND_DIFF_0);

	// Segmento E
	and and10 (SINAL_AND_NOT_DIFF_0, sinal, NOT_DIFF0);
	and and11 (NOT_SINAL_AND_DIFF2, NOT_SINAL, diff[2]);
	and and12 (NOT_DIFF2_AND_DIFF0, NOT_DIFF2, diff[0]);
	or or4 (E, SINAL_AND_NOT_DIFF_0, NOT_SINAL_AND_DIFF3, NOT_SINAL_AND_DIFF2, NOT_DIFF3_AND_DIFF2, NOT_DIFF2_AND_DIFF0);
	
	// Segmento F	
	and and13 (NOT_DIFF3_AND_DIFF1, NOT_DIFF3, diff[1]);
	or or5 (F, SINAL_AND_NOT_DIFF_0, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF1, DIFF2_AND_NOT_DIFF1, NOT_DIFF2_AND_DIFF0);
	
	// Segmento G
	and and14 (SINAL_AND_DIFF1, sinal, diff[1]);
	and and15 (NOT_DIFF2_AND_NOT_DIFF1, NOT_DIFF2, NOT_DIFF1);
	and and16 (NOT_DIFF1_AND_NOT_DIFF0, NOT_DIFF1, NOT_DIFF0);
	
	or or6 (G, SINAL_AND_DIFF1, NOT_SINAL_AND_DIFF3, NOT_DIFF3_AND_DIFF2, NOT_DIFF2_AND_NOT_DIFF1, NOT_DIFF1_AND_NOT_DIFF0);
	
	// Segmento DP
	or or7 (DP, sinal, diff[3], diff[2]);
	
endmodule 